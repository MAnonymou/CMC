module wn1 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp2 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn2 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp3 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn3 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp4 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn4 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp5 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn5 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp6 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn6 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp7 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn7 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp8 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn8 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp9 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn9 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp10 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn10 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp11 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn11 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp12 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn12 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp13 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn13 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp14 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn14 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp15 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn15 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp16 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn16 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp17 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn17 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp18 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn18 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp19 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn19 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp20 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn20 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp21 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn21 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp22 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn22 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp23 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn23 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp24 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn24 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp25 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn25 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp26 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn26 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp27 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn27 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp28 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn28 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp29 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn29 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp30 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn30 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp31 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn31 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp32 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn32 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp33 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn33 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp34 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn34 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp35 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn35 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp36 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn36 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp37 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn37 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp38 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn38 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp39 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn39 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp40 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn40 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp41 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn41 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp42 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn42 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp43 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn43 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp44 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn44 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp45 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn45 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp46 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn46 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp47 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn47 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp48 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn48 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp49 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn49 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp50 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn50 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp51 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn51 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp52 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn52 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp53 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn53 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp54 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn54 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp55 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn55 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp56 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn56 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp57 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn57 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp58 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn58 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp59 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn59 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp60 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn60 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp61 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn61 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp62 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn62 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp63 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn63 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp64 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn64 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp65 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn65 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp66 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn66 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp67 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn67 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp68 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn68 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp69 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn69 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp70 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn70 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp71 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn71 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp72 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn72 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp73 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn73 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp74 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn74 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp75 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn75 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp76 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn76 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp77 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn77 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp78 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn78 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp79 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn79 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp80 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn80 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp81 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn81 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp82 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn82 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp83 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn83 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp84 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn84 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp85 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn85 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp86 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn86 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp87 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn87 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp88 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn88 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp89 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn89 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp90 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn90 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp91 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn91 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp92 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn92 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp93 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn93 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp94 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn94 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp95 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn95 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp96 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn96 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp97 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn97 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp98 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn98 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp99 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn99 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp100 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn100 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp101 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn101 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp102 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn102 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp103 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn103 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp104 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn104 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp105 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn105 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp106 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn106 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp107 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn107 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp108 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn108 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp109 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn109 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp110 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn110 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp111 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn111 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp112 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn112 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp113 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn113 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp114 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn114 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp115 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn115 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp116 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn116 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp117 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn117 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp118 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn118 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp119 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn119 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp120 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn120 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp121 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn121 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp122 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn122 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp123 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn123 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp124 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn124 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp125 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn125 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp126 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn126 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wp127 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= din[7];
end
endmodule

module wn127 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

module wn128 (input [7:0] din, output reg [14:0] dout);
always@(*)
begin
	dout[13:0] <= {din[5:0],din[7:0]};
	dout[14] <= ~ din[7];
end
endmodule

