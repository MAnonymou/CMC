module wn1 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp2 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn2 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp3 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn3 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp4 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn4 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp5 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn5 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp6 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn6 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp7 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn7 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp8 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn8 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp9 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn9 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp10 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn10 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp11 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn11 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp12 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn12 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp13 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn13 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp14 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn14 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp15 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn15 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp16 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn16 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp17 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn17 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp18 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn18 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp19 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn19 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp20 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn20 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp21 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn21 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp22 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn22 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp23 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn23 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp24 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn24 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp25 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn25 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp26 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn26 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp27 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn27 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp28 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn28 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp29 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn29 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp30 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn30 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wp31 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= din[5];
end
endmodule

module wn31 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

module wn32 (input [5:0] din, output reg [10:0] dout);
always@(*)
begin
	dout[9:0] <= {din[3:0],din[5:0]};
	dout[10] <= ~ din[5];
end
endmodule

